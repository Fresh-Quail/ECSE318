module serialAdder(A, B, clear );
parameter N = 6;
input [N-1:0] A, B;
output 